write_pc(32'h10000000);
write_mem(32'h10000000, 32'hFFFC0403);
write_reg(5'd24, 32'h10000104);
write_mem(32'h10000100, 32'hA5000000);
