write_pc(32'h10000000);
write_mem(32'h10000000, 32'h1107C063);
write_reg(5'd15, 32'h00000064);
write_reg(5'd16, 32'h0000000A);