write_pc(32'h10000000);
write_mem(32'h10000000, 32'h10028267);
write_reg(5'h5, 32'h10000000);