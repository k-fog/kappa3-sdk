write_pc(32'h10000000);
write_mem(32'h10000000, 32'h10A48063);
write_reg(5'h9, 32'h0000000A);
write_reg(5'ha, 32'h00000000);