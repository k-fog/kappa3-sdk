write_pc(32'h10000000);
write_mem(32'h10000000, 32'h00942633);
write_reg(5'd8, 32'h0000000A);
write_reg(5'd9, 32'h00000064);
