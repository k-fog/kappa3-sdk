write_pc(32'h10000000);
write_mem(32'h10000000, 32'h10628063);
write_reg(5'h5, 32'h0000000A);
write_reg(5'h6, 32'h0000000A);