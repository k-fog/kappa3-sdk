write_pc(32'h10000000);
write_mem(32'h10000000, 32'h10C5C063);
write_reg(5'd11, 32'h0000000A);
write_reg(5'd12, 32'h00000064);