write_pc(32'h10000000);
write_mem(32'h10000000, 32'h009B0303);
write_reg(5'd22, 32'h100000F8);
write_mem(32'h10000100, 32'h0000A500);
