write_pc(32'h10000000);
write_mem(32'h10000000, 32'hFFCCA483);
write_reg(5'd25, 32'h10000104);
write_mem(32'h10000100, 32'h12345678);
