write_pc(32'h10000000);
write_mem(32'h10000000, 32'h000A8283);
write_reg(5'd21, 32'h10000100);
write_mem(32'h10000100, 32'h000000A5);