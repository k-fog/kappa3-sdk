write_pc(32'h10000000);
write_mem(32'h10000000, 32'h86543117);