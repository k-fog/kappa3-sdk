read_mem(32'h10000100);