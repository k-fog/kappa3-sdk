write_pc(32'h10000000);
write_mem(32'h10000000, 32'h007305B3);
write_reg(5'd6, 32'h0000000A);
write_reg(5'd7, 32'hFFFFFFFD);
