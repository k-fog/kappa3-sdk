write_pc(32'h10000000);
write_mem(32'h10000000, 32'h1149E063);
write_reg(5'd19, 32'hFFFFFFF6);
write_reg(5'd20, 32'h00000064);