write_pc(32'h10000000);
write_mem(32'h10000000, 32'hFFD28513);
write_reg(5'd5, 32'h0000000A);
