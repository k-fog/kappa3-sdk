write_pc(32'h10000000);
write_mem(32'h10000000, 32'h006B8383);
write_reg(5'd23, 32'h100000FC);
write_mem(32'h10000100, 32'h00A50000);
