write_pc(32'h10000000);
write_mem(32'h10000000, 32'hF0E6C0E3);
write_reg(5'd13, 32'hFFFFFFF6);
write_reg(5'd14, 32'h00000064);