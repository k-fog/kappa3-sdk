write_pc(32'h10000000);
write_mem(32'h10000000, 32'hF08380E3);
write_reg(5'h7, 32'h0000000A);
write_reg(5'h8, 32'h0000000A);