write_pc(32'h10000000);
write_mem(32'h10000000, 32'h1128E063);
write_reg(5'd17, 32'h0000000A);
write_reg(5'd18, 32'h00000064);